`include "defines.v"

module brouter_3x3(
    input   `control_w  b0000_ci,
    input   `control_w	b0001_ci,
    input   `control_w	b0010_ci,
    input   `control_w  b0100_ci,
    input   `control_w	b0101_ci,
    input   `control_w	b0110_ci,
    input   `control_w	b1000_ci,
    input   `control_w	b1001_ci,
    input   `control_w	b1010_ci,
    input   `data_w	    b0000_di,
    input   `data_w	    b0001_di,
    input   `data_w 	b0010_di,
    input   `data_w	    b0100_di,
    input   `data_w	    b0101_di,
    input   `data_w	    b0110_di,
    input   `data_w	    b1000_di,
    input   `data_w	    b1001_di,
    input   `data_w     b1010_di,
    input               clk,
    input               rst,
    output  `control_w  b0000_co,
    output  `control_w	b0001_co,
    output  `control_w	b0010_co,
    output  `control_w  b0100_co,
    output  `control_w	b0101_co,
    output  `control_w	b0110_co,
    output  `control_w	b1000_co,
    output  `control_w	b1001_co,
    output  `control_w	b1010_co,
    output  `data_w     b0000_do,
    output  `data_w     b0001_do,
    output  `data_w 	b0010_do,
    output  `data_w     b0100_do,
    output  `data_w     b0101_do,
    output  `data_w     b0110_do,
    output  `data_w     b1000_do,
    output  `data_w     b1001_do,
    output  `data_w     b1010_do,
    output       	    b0000_r,
    output       	    b0001_r,
    output            	b0010_r,
    output       	    b0100_r,
    output       	    b0101_r,
    output       	    b0110_r,
    output       	    b1000_r,
    output       	    b1001_r,
    output       	    b1010_r);

    wire    `control_w  c01, c10, c12, c21, c02, c20,   // Cols
                        c45, c54, c56, c65, c46, c64,
                        c89, c98, ca9, c9a, c8a, ca8,
                        c04, c40, c48, c84, c08, c80,   // Rows
                        c15, c51, c59, c95, c19, c91,
                        c26, c62, c6a, ca6, c2a, ca2;

    wire    `data_w     d01, d10, d12, d21, d02, d20,   // Cols
                        d45, d54, d56, d65, d46, d64,
                        d89, d98, da9, d9a, d8a, da8,
                        d04, d40, d48, d84, d08, d80,   // Rows
                        d15, d51, d59, d95, d19, d91,
                        d26, d62, d6a, da6, d2a, da2;


    brouter #(4'b0000) br0000
                   (.port0_ci(c20),
                    .port0_di(d20),
                    .port0_co(c02),
                    .port0_do(d02),
                    .port1_ci(c10),
                    .port1_di(d10),
                    .port1_co(c01),
                    .port1_do(d01),
                    .port2_ci(c40),
                    .port2_di(d40),
                    .port2_co(c04),
                    .port2_do(d04),
                    .port3_ci(c80),
                    .port3_di(d80),
                    .port3_co(c08),
                    .port3_do(d08),
                    .port4_ci(b0000_ci),
                    .port4_di(b0000_di),
                    .port4_co(b0000_co),
                    .port4_do(b0000_do),
                    .port4_ready(b0000_r),
                    .clk(clk),
                    .rst(rst));
    brouter #(4'b0001) br0001
                   (.port0_ci(c01),
                    .port0_di(d01),
                    .port0_co(c10),
                    .port0_do(d10),
                    .port1_ci(c21),
                    .port1_di(d21),
                    .port1_co(c12),
                    .port1_do(d12),
                    .port2_ci(c51),
                    .port2_di(d51),
                    .port2_co(c15),
                    .port2_do(d15),
                    .port3_ci(c91),
                    .port3_di(d91),
                    .port3_co(c19),
                    .port3_do(d19),
                    .port4_ci(b0001_ci),
                    .port4_di(b0001_di),
                    .port4_co(b0001_co),
                    .port4_do(b0001_do),
                    .port4_ready(b0001_r),
                    .clk(clk),
                    .rst(rst));
    brouter #(4'b0010) br0010 
                   (.port0_ci(c12),
                    .port0_di(d12),
                    .port0_co(c21),
                    .port0_do(d21),
                    .port1_ci(c02),
                    .port1_di(d02),
                    .port1_co(c20),
                    .port1_do(d20),
                    .port2_ci(c62),
                    .port2_di(d62),
                    .port2_co(c26),
                    .port2_do(d26),
                    .port3_ci(ca2),
                    .port3_di(da2),
                    .port3_co(c2a),
                    .port3_do(d2a),
                    .port4_ci(b0010_ci),
                    .port4_di(b0010_di),
                    .port4_co(b0010_co),
                    .port4_do(b0010_do),
                    .port4_ready(b0010_r),
                    .clk(clk),
                    .rst(rst));
    brouter #(4'b0100) br0100
                   (.port0_ci(c64),
                    .port0_di(d64),
                    .port0_co(c46),
                    .port0_do(d46),
                    .port1_ci(c54),
                    .port1_di(d54),
                    .port1_co(c45),
                    .port1_do(d45),
                    .port2_ci(c84),
                    .port2_di(d84),
                    .port2_co(c48),
                    .port2_do(d48),
                    .port3_ci(c04),
                    .port3_di(d04),
                    .port3_co(c40),
                    .port3_do(d40),
                    .port4_ci(b0100_ci),
                    .port4_di(b0100_di),
                    .port4_co(b0100_co),
                    .port4_do(b0100_do),
                    .port4_ready(b0100_r),
                    .clk(clk),
                    .rst(rst));
    brouter #(4'b0101) br0101 
                   (.port0_ci(c45),
                    .port0_di(d45),
                    .port0_co(c54),
                    .port0_do(d54),
                    .port1_ci(c65),
                    .port1_di(d65),
                    .port1_co(c56),
                    .port1_do(d56),
                    .port2_ci(c95),
                    .port2_di(d95),
                    .port2_co(c59),
                    .port2_do(d59),
                    .port3_ci(c15),
                    .port3_di(d15),
                    .port3_co(c51),
                    .port3_do(d51),
                    .port4_ci(b0101_ci),
                    .port4_di(b0101_di),
                    .port4_co(b0101_co),
                    .port4_do(b0101_do),
                    .port4_ready(b0101_r),
                    .clk(clk),
                    .rst(rst));
    brouter #(4'b0110) br0110
                   (.port0_ci(c56),
                    .port0_di(d56),
                    .port0_co(c65),
                    .port0_do(d65),
                    .port1_ci(c46),
                    .port1_di(d46),
                    .port1_co(c64),
                    .port1_do(d64),
                    .port2_ci(ca6),
                    .port2_di(da6),
                    .port2_co(c6a),
                    .port2_do(d6a),
                    .port3_ci(c26),
                    .port3_di(d26),
                    .port3_co(c62),
                    .port3_do(d62),
                    .port4_ci(b0110_ci),
                    .port4_di(b0110_di),
                    .port4_co(b0110_co),
                    .port4_do(b0110_do),
                    .port4_ready(b0110_r),
                    .clk(clk),
                    .rst(rst));
    brouter #(4'b1000) br1000 
                   (.port0_ci(ca8),
                    .port0_di(da8),
                    .port0_co(c8a),
                    .port0_do(d8a),
                    .port1_ci(c98),
                    .port1_di(d98),
                    .port1_co(c89),
                    .port1_do(d89),
                    .port2_ci(c08),
                    .port2_di(d08),
                    .port2_co(c80),
                    .port2_do(d80),
                    .port3_ci(c48),
                    .port3_di(d48),
                    .port3_co(c84),
                    .port3_do(d84),
                    .port4_ci(b1000_ci),
                    .port4_di(b1000_di),
                    .port4_co(b1000_co),
                    .port4_do(b1000_do),
                    .port4_ready(b1000_r),
                    .clk(clk),
                    .rst(rst));
    brouter #(4'b1001) br1001 
                   (.port0_ci(c89),
                    .port0_di(d89),
                    .port0_co(c98),
                    .port0_do(d98),
                    .port1_ci(ca9),
                    .port1_di(da9),
                    .port1_co(c9a),
                    .port1_do(d9a),
                    .port2_ci(c19),
                    .port2_di(d19),
                    .port2_co(c91),
                    .port2_do(d91),
                    .port3_ci(c59),
                    .port3_di(d59),
                    .port3_co(c95),
                    .port3_do(d95),
                    .port4_ci(b1001_ci),
                    .port4_di(b1001_di),
                    .port4_co(b1001_co),
                    .port4_do(b1001_do),
                    .port4_ready(b1001_r),
                    .clk(clk),
                    .rst(rst));
    brouter #(4'b1010) br1010 
                   (.port0_ci(c9a),
                    .port0_di(d9a),
                    .port0_co(ca9),
                    .port0_do(da9),
                    .port1_ci(c8a),
                    .port1_di(d8a),
                    .port1_co(ca8),
                    .port1_do(da8),
                    .port2_ci(c2a),
                    .port2_di(d2a),
                    .port2_co(ca2),
                    .port2_do(da2),
                    .port3_ci(c6a),
                    .port3_di(d6a),
                    .port3_co(ca6),
                    .port3_do(da6),
                    .port4_ci(b1010_ci),
                    .port4_di(b1010_di),
                    .port4_co(b1010_co),
                    .port4_do(b1010_do),
                    .port4_ready(b1010_r),
                    .clk(clk),
                    .rst(rst));

endmodule
