parameter DIM = 4;           // size in one dimension
parameter ADDRBITS2 = 4;     // bits in two dimensions of address
parameter ADDRBITS = 2;      // bits in one dimension of address
parameter HOPBITS = 8;       // bits for hop-count
parameter LINKWIDTH = 134;   // data bits (128 bits) + header bits (2 bits for type, 1 for length, 3 for flitNr)
